library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package prog_mem is
    type RAM_Array is array (0 to 32767) of std_logic_vector(7 downto 0);
    constant RAM_INIT : RAM_Array := (
        -- LEA R6, start of .TEXT
        16#000# => X"B6", -- opcode LEA R6
        16#001# => X"EE", -- LSB address
        16#002# => X"00", -- MSB address

        -- SECTION .TEXT
        16#0EE# => X"63", -- 238
        16#0EF# => X"04", -- 239
        16#0F0# => X"83", -- 240
        16#0F1# => X"F2", -- 241
        16#0F2# => X"FF", -- 242
        16#0F3# => X"83", -- 243
        16#0F4# => X"F3", -- 244
        16#0F5# => X"FF", -- 245
        16#0F6# => X"71", -- 246
        16#0F7# => X"F4", -- 247
        16#0F8# => X"FF", -- 248
        16#0F9# => X"21", -- 249
        16#0FA# => X"05", -- 250
        16#0FB# => X"96", -- 251
        16#0FC# => X"F6", -- 252
        16#0FD# => X"00", -- 253
        16#0FE# => X"B6", -- 254
        16#0FF# => X"0C", -- 255
        16#100# => X"01", -- 256
        16#101# => X"71", -- 257
        16#102# => X"F4", -- 258
        16#103# => X"FF", -- 259
        16#104# => X"21", -- 260
        16#105# => X"01", -- 261
        16#106# => X"96", -- 262
        16#107# => X"01", -- 263
        16#108# => X"01", -- 264
        16#109# => X"B6", -- 265
        16#10A# => X"1C", -- 266
        16#10B# => X"01", -- 267
        16#10C# => X"63", -- 268
        16#10D# => X"00", -- 269
        16#10E# => X"83", -- 270
        16#10F# => X"F3", -- 271
        16#110# => X"FF", -- 272
        16#111# => X"71", -- 273
        16#112# => X"F4", -- 274
        16#113# => X"FF", -- 275
        16#114# => X"21", -- 276
        16#115# => X"03", -- 277
        16#116# => X"96", -- 278
        16#117# => X"11", -- 279
        16#118# => X"01", -- 280
        16#119# => X"B6", -- 281
        16#11A# => X"01", -- 282
        16#11B# => X"01", -- 283
        16#11C# => X"63", -- 284
        16#11D# => X"04", -- 285
        16#11E# => X"83", -- 286
        16#11F# => X"F3", -- 287
        16#120# => X"FF", -- 288
        16#121# => X"71", -- 289
        16#122# => X"F4", -- 290
        16#123# => X"FF", -- 291
        16#124# => X"21", -- 292
        16#125# => X"07", -- 293
        16#126# => X"96", -- 294
        16#127# => X"21", -- 295
        16#128# => X"01", -- 296
        16#129# => X"B6", -- 297
        16#12A# => X"F6", -- 298
        16#12B# => X"00", -- 299
        16#12C# => X"B6", -- 300
        16#12D# => X"2C", -- 301
        16#12E# => X"01", -- 302

        others => (others => '0')
    );
end package;
